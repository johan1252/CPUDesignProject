--Testbench used to test the CPU_Bus
LIBRARY ieee;
USE ieee.std_logic_1164.all; 

Entity CPU_Bus_tb is
end

Architecture CPU_Bus_tb_arch of CPU_Bus_tb is
signal 