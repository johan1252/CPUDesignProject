-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Tue Jan 26 13:07:55 2016"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Bus IS 
	PORT
	(

	);
END Bus;

ARCHITECTURE bdf_type OF Bus IS 

COMPONENT lpm_encoder
	PORT(eq0 : IN STD_LOGIC;
		 eq1 : IN STD_LOGIC;
		 eq2 : IN STD_LOGIC;
		 eq3 : IN STD_LOGIC;
		 eq4 : IN STD_LOGIC;
		 eq5 : IN STD_LOGIC;
		 eq6 : IN STD_LOGIC;
		 eq7 : IN STD_LOGIC;
		 eq8 : IN STD_LOGIC;
		 eq9 : IN STD_LOGIC;
		 eq10 : IN STD_LOGIC;
		 eq11 : IN STD_LOGIC;
		 eq12 : IN STD_LOGIC;
		 eq13 : IN STD_LOGIC;
		 eq14 : IN STD_LOGIC;
		 eq15 : IN STD_LOGIC;
		 eq16 : IN STD_LOGIC;
		 eq17 : IN STD_LOGIC;
		 eq18 : IN STD_LOGIC;
		 eq19 : IN STD_LOGIC;
		 eq20 : IN STD_LOGIC;
		 eq21 : IN STD_LOGIC;
		 eq22 : IN STD_LOGIC;
		 eq23 : IN STD_LOGIC;
		 eq24 : IN STD_LOGIC;
		 eq25 : IN STD_LOGIC;
		 eq26 : IN STD_LOGIC;
		 eq27 : IN STD_LOGIC;
		 eq28 : IN STD_LOGIC;
		 eq29 : IN STD_LOGIC;
		 eq30 : IN STD_LOGIC;
		 eq31 : IN STD_LOGIC;
		 data : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_mux0
	PORT(data0x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data10x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data11x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data12x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data13x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data14x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data15x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data16x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data17x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data18x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data19x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data20x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data21x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data22x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data23x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data24x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data25x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data26x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data27x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data28x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data29x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data30x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data31x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data4x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data5x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data6x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data7x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data8x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 data9x : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mdr_unit
	PORT(ENABLE : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;
		 READ_MUX : IN STD_LOGIC;
		 MDR_IN_0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MDR_IN_1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MDR_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT reg32
	PORT(ENABLE : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;
		 D_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	BusMuxIn-Hi :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-In_Port :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-Lo :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-MDR :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR0 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR1 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR10 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR11 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR12 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR13 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR14 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR15 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR16 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR17 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR18 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR19 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR2 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR20 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR21 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR22 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR23 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR24 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR25 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR26 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR27 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR28 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR29 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR3 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR30 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR31 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR4 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR5 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR6 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR7 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR8 :  STD_LOGIC;
SIGNAL	BusMuxIn-MDR9 :  STD_LOGIC;
SIGNAL	BusMuxIn-PC :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-R0 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-R10 :  STD_LOGIC;
SIGNAL	BusMuxIn-R100 :  STD_LOGIC;
SIGNAL	BusMuxIn-R101 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1010 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1011 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1012 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1013 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1014 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1015 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1016 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1017 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1018 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1019 :  STD_LOGIC;
SIGNAL	BusMuxIn-R102 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1020 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1021 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1022 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1023 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1024 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1025 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1026 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1027 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1028 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1029 :  STD_LOGIC;
SIGNAL	BusMuxIn-R103 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1030 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1031 :  STD_LOGIC;
SIGNAL	BusMuxIn-R104 :  STD_LOGIC;
SIGNAL	BusMuxIn-R105 :  STD_LOGIC;
SIGNAL	BusMuxIn-R106 :  STD_LOGIC;
SIGNAL	BusMuxIn-R107 :  STD_LOGIC;
SIGNAL	BusMuxIn-R108 :  STD_LOGIC;
SIGNAL	BusMuxIn-R109 :  STD_LOGIC;
SIGNAL	BusMuxIn-R11 :  STD_LOGIC;
SIGNAL	BusMuxIn-R110 :  STD_LOGIC;
SIGNAL	BusMuxIn-R111 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1110 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1111 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1112 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1113 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1114 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1115 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1116 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1117 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1118 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1119 :  STD_LOGIC;
SIGNAL	BusMuxIn-R112 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1120 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1121 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1122 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1123 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1124 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1125 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1126 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1127 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1128 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1129 :  STD_LOGIC;
SIGNAL	BusMuxIn-R113 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1130 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1131 :  STD_LOGIC;
SIGNAL	BusMuxIn-R114 :  STD_LOGIC;
SIGNAL	BusMuxIn-R115 :  STD_LOGIC;
SIGNAL	BusMuxIn-R116 :  STD_LOGIC;
SIGNAL	BusMuxIn-R117 :  STD_LOGIC;
SIGNAL	BusMuxIn-R118 :  STD_LOGIC;
SIGNAL	BusMuxIn-R119 :  STD_LOGIC;
SIGNAL	BusMuxIn-R12 :  STD_LOGIC;
SIGNAL	BusMuxIn-R120 :  STD_LOGIC;
SIGNAL	BusMuxIn-R121 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1210 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1211 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1212 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1213 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1214 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1215 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1216 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1217 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1218 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1219 :  STD_LOGIC;
SIGNAL	BusMuxIn-R122 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1220 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1221 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1222 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1223 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1224 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1225 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1226 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1227 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1228 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1229 :  STD_LOGIC;
SIGNAL	BusMuxIn-R123 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1230 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1231 :  STD_LOGIC;
SIGNAL	BusMuxIn-R124 :  STD_LOGIC;
SIGNAL	BusMuxIn-R125 :  STD_LOGIC;
SIGNAL	BusMuxIn-R126 :  STD_LOGIC;
SIGNAL	BusMuxIn-R127 :  STD_LOGIC;
SIGNAL	BusMuxIn-R128 :  STD_LOGIC;
SIGNAL	BusMuxIn-R129 :  STD_LOGIC;
SIGNAL	BusMuxIn-R13 :  STD_LOGIC;
SIGNAL	BusMuxIn-R130 :  STD_LOGIC;
SIGNAL	BusMuxIn-R131 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1310 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1311 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1312 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1313 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1314 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1315 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1316 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1317 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1318 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1319 :  STD_LOGIC;
SIGNAL	BusMuxIn-R132 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1320 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1321 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1322 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1323 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1324 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1325 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1326 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1327 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1328 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1329 :  STD_LOGIC;
SIGNAL	BusMuxIn-R133 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1330 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1331 :  STD_LOGIC;
SIGNAL	BusMuxIn-R134 :  STD_LOGIC;
SIGNAL	BusMuxIn-R135 :  STD_LOGIC;
SIGNAL	BusMuxIn-R136 :  STD_LOGIC;
SIGNAL	BusMuxIn-R137 :  STD_LOGIC;
SIGNAL	BusMuxIn-R138 :  STD_LOGIC;
SIGNAL	BusMuxIn-R139 :  STD_LOGIC;
SIGNAL	BusMuxIn-R14 :  STD_LOGIC;
SIGNAL	BusMuxIn-R140 :  STD_LOGIC;
SIGNAL	BusMuxIn-R141 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1410 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1411 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1412 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1413 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1414 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1415 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1416 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1417 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1418 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1419 :  STD_LOGIC;
SIGNAL	BusMuxIn-R142 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1420 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1421 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1422 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1423 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1424 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1425 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1426 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1427 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1428 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1429 :  STD_LOGIC;
SIGNAL	BusMuxIn-R143 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1430 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1431 :  STD_LOGIC;
SIGNAL	BusMuxIn-R144 :  STD_LOGIC;
SIGNAL	BusMuxIn-R145 :  STD_LOGIC;
SIGNAL	BusMuxIn-R146 :  STD_LOGIC;
SIGNAL	BusMuxIn-R147 :  STD_LOGIC;
SIGNAL	BusMuxIn-R148 :  STD_LOGIC;
SIGNAL	BusMuxIn-R149 :  STD_LOGIC;
SIGNAL	BusMuxIn-R15 :  STD_LOGIC;
SIGNAL	BusMuxIn-R150 :  STD_LOGIC;
SIGNAL	BusMuxIn-R151 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1510 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1511 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1512 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1513 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1514 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1515 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1516 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1517 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1518 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1519 :  STD_LOGIC;
SIGNAL	BusMuxIn-R152 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1520 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1521 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1522 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1523 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1524 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1525 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1526 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1527 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1528 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1529 :  STD_LOGIC;
SIGNAL	BusMuxIn-R153 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1530 :  STD_LOGIC;
SIGNAL	BusMuxIn-R1531 :  STD_LOGIC;
SIGNAL	BusMuxIn-R154 :  STD_LOGIC;
SIGNAL	BusMuxIn-R155 :  STD_LOGIC;
SIGNAL	BusMuxIn-R156 :  STD_LOGIC;
SIGNAL	BusMuxIn-R157 :  STD_LOGIC;
SIGNAL	BusMuxIn-R158 :  STD_LOGIC;
SIGNAL	BusMuxIn-R159 :  STD_LOGIC;
SIGNAL	BusMuxIn-R16 :  STD_LOGIC;
SIGNAL	BusMuxIn-R17 :  STD_LOGIC;
SIGNAL	BusMuxIn-R18 :  STD_LOGIC;
SIGNAL	BusMuxIn-R19 :  STD_LOGIC;
SIGNAL	BusMuxIn-R2 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-R3 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-R4 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-R5 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-R6 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-R7 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-R8 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-R9 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-ZHi :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn-ZLo :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxIn_Csign :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	BusMuxOut :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	Cout :  STD_LOGIC;
SIGNAL	HIout :  STD_LOGIC;
SIGNAL	In_Portout :  STD_LOGIC;
SIGNAL	LOout :  STD_LOGIC;
SIGNAL	Mdatain :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	MDRout :  STD_LOGIC;
SIGNAL	muxSelect :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL	PCout :  STD_LOGIC;
SIGNAL	R0out :  STD_LOGIC;
SIGNAL	R10out :  STD_LOGIC;
SIGNAL	R11out :  STD_LOGIC;
SIGNAL	R12out :  STD_LOGIC;
SIGNAL	R13out :  STD_LOGIC;
SIGNAL	R14out :  STD_LOGIC;
SIGNAL	R15out :  STD_LOGIC;
SIGNAL	R1out :  STD_LOGIC;
SIGNAL	R2out :  STD_LOGIC;
SIGNAL	R3out :  STD_LOGIC;
SIGNAL	R4out :  STD_LOGIC;
SIGNAL	R5out :  STD_LOGIC;
SIGNAL	R6out :  STD_LOGIC;
SIGNAL	R7out :  STD_LOGIC;
SIGNAL	R8out :  STD_LOGIC;
SIGNAL	R9out :  STD_LOGIC;
SIGNAL	Zhighout :  STD_LOGIC;
SIGNAL	Zlowout :  STD_LOGIC;

SIGNAL	GDFX_TEMP_SIGNAL_5 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_14 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_4 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_13 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_3 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_12 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_2 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_11 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_1 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_10 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_0 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_9 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_6 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_8 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_7 :  STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN 

GDFX_TEMP_SIGNAL_5 <= (BusMuxIn-R1531 & BusMuxIn-R1530 & BusMuxIn-R1529 & BusMuxIn-R1528 & BusMuxIn-R1527 & BusMuxIn-R1526 & BusMuxIn-R1525 & BusMuxIn-R1524 & BusMuxIn-R1523 & BusMuxIn-R1522 & BusMuxIn-R1521 & BusMuxIn-R1520 & BusMuxIn-R1519 & BusMuxIn-R1518 & BusMuxIn-R1517 & BusMuxIn-R1516 & BusMuxIn-R1515 & BusMuxIn-R1514 & BusMuxIn-R1513 & BusMuxIn-R1512 & BusMuxIn-R1511 & BusMuxIn-R1510 & BusMuxIn-R159 & BusMuxIn-R158 & BusMuxIn-R157 & BusMuxIn-R156 & BusMuxIn-R155 & BusMuxIn-R154 & BusMuxIn-R153 & BusMuxIn-R152 & BusMuxIn-R151 & BusMuxIn-R150);
BusMuxIn-R1531 <= GDFX_TEMP_SIGNAL_14(31);
BusMuxIn-R1530 <= GDFX_TEMP_SIGNAL_14(30);
BusMuxIn-R1529 <= GDFX_TEMP_SIGNAL_14(29);
BusMuxIn-R1528 <= GDFX_TEMP_SIGNAL_14(28);
BusMuxIn-R1527 <= GDFX_TEMP_SIGNAL_14(27);
BusMuxIn-R1526 <= GDFX_TEMP_SIGNAL_14(26);
BusMuxIn-R1525 <= GDFX_TEMP_SIGNAL_14(25);
BusMuxIn-R1524 <= GDFX_TEMP_SIGNAL_14(24);
BusMuxIn-R1523 <= GDFX_TEMP_SIGNAL_14(23);
BusMuxIn-R1522 <= GDFX_TEMP_SIGNAL_14(22);
BusMuxIn-R1521 <= GDFX_TEMP_SIGNAL_14(21);
BusMuxIn-R1520 <= GDFX_TEMP_SIGNAL_14(20);
BusMuxIn-R1519 <= GDFX_TEMP_SIGNAL_14(19);
BusMuxIn-R1518 <= GDFX_TEMP_SIGNAL_14(18);
BusMuxIn-R1517 <= GDFX_TEMP_SIGNAL_14(17);
BusMuxIn-R1516 <= GDFX_TEMP_SIGNAL_14(16);
BusMuxIn-R1515 <= GDFX_TEMP_SIGNAL_14(15);
BusMuxIn-R1514 <= GDFX_TEMP_SIGNAL_14(14);
BusMuxIn-R1513 <= GDFX_TEMP_SIGNAL_14(13);
BusMuxIn-R1512 <= GDFX_TEMP_SIGNAL_14(12);
BusMuxIn-R1511 <= GDFX_TEMP_SIGNAL_14(11);
BusMuxIn-R1510 <= GDFX_TEMP_SIGNAL_14(10);
BusMuxIn-R159 <= GDFX_TEMP_SIGNAL_14(9);
BusMuxIn-R158 <= GDFX_TEMP_SIGNAL_14(8);
BusMuxIn-R157 <= GDFX_TEMP_SIGNAL_14(7);
BusMuxIn-R156 <= GDFX_TEMP_SIGNAL_14(6);
BusMuxIn-R155 <= GDFX_TEMP_SIGNAL_14(5);
BusMuxIn-R154 <= GDFX_TEMP_SIGNAL_14(4);
BusMuxIn-R153 <= GDFX_TEMP_SIGNAL_14(3);
BusMuxIn-R152 <= GDFX_TEMP_SIGNAL_14(2);
BusMuxIn-R151 <= GDFX_TEMP_SIGNAL_14(1);
BusMuxIn-R150 <= GDFX_TEMP_SIGNAL_14(0);

GDFX_TEMP_SIGNAL_4 <= (BusMuxIn-R1431 & BusMuxIn-R1430 & BusMuxIn-R1429 & BusMuxIn-R1428 & BusMuxIn-R1427 & BusMuxIn-R1426 & BusMuxIn-R1425 & BusMuxIn-R1424 & BusMuxIn-R1423 & BusMuxIn-R1422 & BusMuxIn-R1421 & BusMuxIn-R1420 & BusMuxIn-R1419 & BusMuxIn-R1418 & BusMuxIn-R1417 & BusMuxIn-R1416 & BusMuxIn-R1415 & BusMuxIn-R1414 & BusMuxIn-R1413 & BusMuxIn-R1412 & BusMuxIn-R1411 & BusMuxIn-R1410 & BusMuxIn-R149 & BusMuxIn-R148 & BusMuxIn-R147 & BusMuxIn-R146 & BusMuxIn-R145 & BusMuxIn-R144 & BusMuxIn-R143 & BusMuxIn-R142 & BusMuxIn-R141 & BusMuxIn-R140);
BusMuxIn-R1431 <= GDFX_TEMP_SIGNAL_13(31);
BusMuxIn-R1430 <= GDFX_TEMP_SIGNAL_13(30);
BusMuxIn-R1429 <= GDFX_TEMP_SIGNAL_13(29);
BusMuxIn-R1428 <= GDFX_TEMP_SIGNAL_13(28);
BusMuxIn-R1427 <= GDFX_TEMP_SIGNAL_13(27);
BusMuxIn-R1426 <= GDFX_TEMP_SIGNAL_13(26);
BusMuxIn-R1425 <= GDFX_TEMP_SIGNAL_13(25);
BusMuxIn-R1424 <= GDFX_TEMP_SIGNAL_13(24);
BusMuxIn-R1423 <= GDFX_TEMP_SIGNAL_13(23);
BusMuxIn-R1422 <= GDFX_TEMP_SIGNAL_13(22);
BusMuxIn-R1421 <= GDFX_TEMP_SIGNAL_13(21);
BusMuxIn-R1420 <= GDFX_TEMP_SIGNAL_13(20);
BusMuxIn-R1419 <= GDFX_TEMP_SIGNAL_13(19);
BusMuxIn-R1418 <= GDFX_TEMP_SIGNAL_13(18);
BusMuxIn-R1417 <= GDFX_TEMP_SIGNAL_13(17);
BusMuxIn-R1416 <= GDFX_TEMP_SIGNAL_13(16);
BusMuxIn-R1415 <= GDFX_TEMP_SIGNAL_13(15);
BusMuxIn-R1414 <= GDFX_TEMP_SIGNAL_13(14);
BusMuxIn-R1413 <= GDFX_TEMP_SIGNAL_13(13);
BusMuxIn-R1412 <= GDFX_TEMP_SIGNAL_13(12);
BusMuxIn-R1411 <= GDFX_TEMP_SIGNAL_13(11);
BusMuxIn-R1410 <= GDFX_TEMP_SIGNAL_13(10);
BusMuxIn-R149 <= GDFX_TEMP_SIGNAL_13(9);
BusMuxIn-R148 <= GDFX_TEMP_SIGNAL_13(8);
BusMuxIn-R147 <= GDFX_TEMP_SIGNAL_13(7);
BusMuxIn-R146 <= GDFX_TEMP_SIGNAL_13(6);
BusMuxIn-R145 <= GDFX_TEMP_SIGNAL_13(5);
BusMuxIn-R144 <= GDFX_TEMP_SIGNAL_13(4);
BusMuxIn-R143 <= GDFX_TEMP_SIGNAL_13(3);
BusMuxIn-R142 <= GDFX_TEMP_SIGNAL_13(2);
BusMuxIn-R141 <= GDFX_TEMP_SIGNAL_13(1);
BusMuxIn-R140 <= GDFX_TEMP_SIGNAL_13(0);

GDFX_TEMP_SIGNAL_3 <= (BusMuxIn-R1331 & BusMuxIn-R1330 & BusMuxIn-R1329 & BusMuxIn-R1328 & BusMuxIn-R1327 & BusMuxIn-R1326 & BusMuxIn-R1325 & BusMuxIn-R1324 & BusMuxIn-R1323 & BusMuxIn-R1322 & BusMuxIn-R1321 & BusMuxIn-R1320 & BusMuxIn-R1319 & BusMuxIn-R1318 & BusMuxIn-R1317 & BusMuxIn-R1316 & BusMuxIn-R1315 & BusMuxIn-R1314 & BusMuxIn-R1313 & BusMuxIn-R1312 & BusMuxIn-R1311 & BusMuxIn-R1310 & BusMuxIn-R139 & BusMuxIn-R138 & BusMuxIn-R137 & BusMuxIn-R136 & BusMuxIn-R135 & BusMuxIn-R134 & BusMuxIn-R133 & BusMuxIn-R132 & BusMuxIn-R131 & BusMuxIn-R130);
BusMuxIn-R1331 <= GDFX_TEMP_SIGNAL_12(31);
BusMuxIn-R1330 <= GDFX_TEMP_SIGNAL_12(30);
BusMuxIn-R1329 <= GDFX_TEMP_SIGNAL_12(29);
BusMuxIn-R1328 <= GDFX_TEMP_SIGNAL_12(28);
BusMuxIn-R1327 <= GDFX_TEMP_SIGNAL_12(27);
BusMuxIn-R1326 <= GDFX_TEMP_SIGNAL_12(26);
BusMuxIn-R1325 <= GDFX_TEMP_SIGNAL_12(25);
BusMuxIn-R1324 <= GDFX_TEMP_SIGNAL_12(24);
BusMuxIn-R1323 <= GDFX_TEMP_SIGNAL_12(23);
BusMuxIn-R1322 <= GDFX_TEMP_SIGNAL_12(22);
BusMuxIn-R1321 <= GDFX_TEMP_SIGNAL_12(21);
BusMuxIn-R1320 <= GDFX_TEMP_SIGNAL_12(20);
BusMuxIn-R1319 <= GDFX_TEMP_SIGNAL_12(19);
BusMuxIn-R1318 <= GDFX_TEMP_SIGNAL_12(18);
BusMuxIn-R1317 <= GDFX_TEMP_SIGNAL_12(17);
BusMuxIn-R1316 <= GDFX_TEMP_SIGNAL_12(16);
BusMuxIn-R1315 <= GDFX_TEMP_SIGNAL_12(15);
BusMuxIn-R1314 <= GDFX_TEMP_SIGNAL_12(14);
BusMuxIn-R1313 <= GDFX_TEMP_SIGNAL_12(13);
BusMuxIn-R1312 <= GDFX_TEMP_SIGNAL_12(12);
BusMuxIn-R1311 <= GDFX_TEMP_SIGNAL_12(11);
BusMuxIn-R1310 <= GDFX_TEMP_SIGNAL_12(10);
BusMuxIn-R139 <= GDFX_TEMP_SIGNAL_12(9);
BusMuxIn-R138 <= GDFX_TEMP_SIGNAL_12(8);
BusMuxIn-R137 <= GDFX_TEMP_SIGNAL_12(7);
BusMuxIn-R136 <= GDFX_TEMP_SIGNAL_12(6);
BusMuxIn-R135 <= GDFX_TEMP_SIGNAL_12(5);
BusMuxIn-R134 <= GDFX_TEMP_SIGNAL_12(4);
BusMuxIn-R133 <= GDFX_TEMP_SIGNAL_12(3);
BusMuxIn-R132 <= GDFX_TEMP_SIGNAL_12(2);
BusMuxIn-R131 <= GDFX_TEMP_SIGNAL_12(1);
BusMuxIn-R130 <= GDFX_TEMP_SIGNAL_12(0);

GDFX_TEMP_SIGNAL_2 <= (BusMuxIn-R1231 & BusMuxIn-R1230 & BusMuxIn-R1229 & BusMuxIn-R1228 & BusMuxIn-R1227 & BusMuxIn-R1226 & BusMuxIn-R1225 & BusMuxIn-R1224 & BusMuxIn-R1223 & BusMuxIn-R1222 & BusMuxIn-R1221 & BusMuxIn-R1220 & BusMuxIn-R1219 & BusMuxIn-R1218 & BusMuxIn-R1217 & BusMuxIn-R1216 & BusMuxIn-R1215 & BusMuxIn-R1214 & BusMuxIn-R1213 & BusMuxIn-R1212 & BusMuxIn-R1211 & BusMuxIn-R1210 & BusMuxIn-R129 & BusMuxIn-R128 & BusMuxIn-R127 & BusMuxIn-R126 & BusMuxIn-R125 & BusMuxIn-R124 & BusMuxIn-R123 & BusMuxIn-R122 & BusMuxIn-R121 & BusMuxIn-R120);
BusMuxIn-R1231 <= GDFX_TEMP_SIGNAL_11(31);
BusMuxIn-R1230 <= GDFX_TEMP_SIGNAL_11(30);
BusMuxIn-R1229 <= GDFX_TEMP_SIGNAL_11(29);
BusMuxIn-R1228 <= GDFX_TEMP_SIGNAL_11(28);
BusMuxIn-R1227 <= GDFX_TEMP_SIGNAL_11(27);
BusMuxIn-R1226 <= GDFX_TEMP_SIGNAL_11(26);
BusMuxIn-R1225 <= GDFX_TEMP_SIGNAL_11(25);
BusMuxIn-R1224 <= GDFX_TEMP_SIGNAL_11(24);
BusMuxIn-R1223 <= GDFX_TEMP_SIGNAL_11(23);
BusMuxIn-R1222 <= GDFX_TEMP_SIGNAL_11(22);
BusMuxIn-R1221 <= GDFX_TEMP_SIGNAL_11(21);
BusMuxIn-R1220 <= GDFX_TEMP_SIGNAL_11(20);
BusMuxIn-R1219 <= GDFX_TEMP_SIGNAL_11(19);
BusMuxIn-R1218 <= GDFX_TEMP_SIGNAL_11(18);
BusMuxIn-R1217 <= GDFX_TEMP_SIGNAL_11(17);
BusMuxIn-R1216 <= GDFX_TEMP_SIGNAL_11(16);
BusMuxIn-R1215 <= GDFX_TEMP_SIGNAL_11(15);
BusMuxIn-R1214 <= GDFX_TEMP_SIGNAL_11(14);
BusMuxIn-R1213 <= GDFX_TEMP_SIGNAL_11(13);
BusMuxIn-R1212 <= GDFX_TEMP_SIGNAL_11(12);
BusMuxIn-R1211 <= GDFX_TEMP_SIGNAL_11(11);
BusMuxIn-R1210 <= GDFX_TEMP_SIGNAL_11(10);
BusMuxIn-R129 <= GDFX_TEMP_SIGNAL_11(9);
BusMuxIn-R128 <= GDFX_TEMP_SIGNAL_11(8);
BusMuxIn-R127 <= GDFX_TEMP_SIGNAL_11(7);
BusMuxIn-R126 <= GDFX_TEMP_SIGNAL_11(6);
BusMuxIn-R125 <= GDFX_TEMP_SIGNAL_11(5);
BusMuxIn-R124 <= GDFX_TEMP_SIGNAL_11(4);
BusMuxIn-R123 <= GDFX_TEMP_SIGNAL_11(3);
BusMuxIn-R122 <= GDFX_TEMP_SIGNAL_11(2);
BusMuxIn-R121 <= GDFX_TEMP_SIGNAL_11(1);
BusMuxIn-R120 <= GDFX_TEMP_SIGNAL_11(0);

GDFX_TEMP_SIGNAL_1 <= (BusMuxIn-R1131 & BusMuxIn-R1130 & BusMuxIn-R1129 & BusMuxIn-R1128 & BusMuxIn-R1127 & BusMuxIn-R1126 & BusMuxIn-R1125 & BusMuxIn-R1124 & BusMuxIn-R1123 & BusMuxIn-R1122 & BusMuxIn-R1121 & BusMuxIn-R1120 & BusMuxIn-R1119 & BusMuxIn-R1118 & BusMuxIn-R1117 & BusMuxIn-R1116 & BusMuxIn-R1115 & BusMuxIn-R1114 & BusMuxIn-R1113 & BusMuxIn-R1112 & BusMuxIn-R1111 & BusMuxIn-R1110 & BusMuxIn-R119 & BusMuxIn-R118 & BusMuxIn-R117 & BusMuxIn-R116 & BusMuxIn-R115 & BusMuxIn-R114 & BusMuxIn-R113 & BusMuxIn-R112 & BusMuxIn-R111 & BusMuxIn-R110);
BusMuxIn-R1131 <= GDFX_TEMP_SIGNAL_10(31);
BusMuxIn-R1130 <= GDFX_TEMP_SIGNAL_10(30);
BusMuxIn-R1129 <= GDFX_TEMP_SIGNAL_10(29);
BusMuxIn-R1128 <= GDFX_TEMP_SIGNAL_10(28);
BusMuxIn-R1127 <= GDFX_TEMP_SIGNAL_10(27);
BusMuxIn-R1126 <= GDFX_TEMP_SIGNAL_10(26);
BusMuxIn-R1125 <= GDFX_TEMP_SIGNAL_10(25);
BusMuxIn-R1124 <= GDFX_TEMP_SIGNAL_10(24);
BusMuxIn-R1123 <= GDFX_TEMP_SIGNAL_10(23);
BusMuxIn-R1122 <= GDFX_TEMP_SIGNAL_10(22);
BusMuxIn-R1121 <= GDFX_TEMP_SIGNAL_10(21);
BusMuxIn-R1120 <= GDFX_TEMP_SIGNAL_10(20);
BusMuxIn-R1119 <= GDFX_TEMP_SIGNAL_10(19);
BusMuxIn-R1118 <= GDFX_TEMP_SIGNAL_10(18);
BusMuxIn-R1117 <= GDFX_TEMP_SIGNAL_10(17);
BusMuxIn-R1116 <= GDFX_TEMP_SIGNAL_10(16);
BusMuxIn-R1115 <= GDFX_TEMP_SIGNAL_10(15);
BusMuxIn-R1114 <= GDFX_TEMP_SIGNAL_10(14);
BusMuxIn-R1113 <= GDFX_TEMP_SIGNAL_10(13);
BusMuxIn-R1112 <= GDFX_TEMP_SIGNAL_10(12);
BusMuxIn-R1111 <= GDFX_TEMP_SIGNAL_10(11);
BusMuxIn-R1110 <= GDFX_TEMP_SIGNAL_10(10);
BusMuxIn-R119 <= GDFX_TEMP_SIGNAL_10(9);
BusMuxIn-R118 <= GDFX_TEMP_SIGNAL_10(8);
BusMuxIn-R117 <= GDFX_TEMP_SIGNAL_10(7);
BusMuxIn-R116 <= GDFX_TEMP_SIGNAL_10(6);
BusMuxIn-R115 <= GDFX_TEMP_SIGNAL_10(5);
BusMuxIn-R114 <= GDFX_TEMP_SIGNAL_10(4);
BusMuxIn-R113 <= GDFX_TEMP_SIGNAL_10(3);
BusMuxIn-R112 <= GDFX_TEMP_SIGNAL_10(2);
BusMuxIn-R111 <= GDFX_TEMP_SIGNAL_10(1);
BusMuxIn-R110 <= GDFX_TEMP_SIGNAL_10(0);

GDFX_TEMP_SIGNAL_0 <= (BusMuxIn-R1031 & BusMuxIn-R1030 & BusMuxIn-R1029 & BusMuxIn-R1028 & BusMuxIn-R1027 & BusMuxIn-R1026 & BusMuxIn-R1025 & BusMuxIn-R1024 & BusMuxIn-R1023 & BusMuxIn-R1022 & BusMuxIn-R1021 & BusMuxIn-R1020 & BusMuxIn-R1019 & BusMuxIn-R1018 & BusMuxIn-R1017 & BusMuxIn-R1016 & BusMuxIn-R1015 & BusMuxIn-R1014 & BusMuxIn-R1013 & BusMuxIn-R1012 & BusMuxIn-R1011 & BusMuxIn-R1010 & BusMuxIn-R109 & BusMuxIn-R108 & BusMuxIn-R107 & BusMuxIn-R106 & BusMuxIn-R105 & BusMuxIn-R104 & BusMuxIn-R103 & BusMuxIn-R102 & BusMuxIn-R101 & BusMuxIn-R100);
BusMuxIn-R1031 <= GDFX_TEMP_SIGNAL_9(31);
BusMuxIn-R1030 <= GDFX_TEMP_SIGNAL_9(30);
BusMuxIn-R1029 <= GDFX_TEMP_SIGNAL_9(29);
BusMuxIn-R1028 <= GDFX_TEMP_SIGNAL_9(28);
BusMuxIn-R1027 <= GDFX_TEMP_SIGNAL_9(27);
BusMuxIn-R1026 <= GDFX_TEMP_SIGNAL_9(26);
BusMuxIn-R1025 <= GDFX_TEMP_SIGNAL_9(25);
BusMuxIn-R1024 <= GDFX_TEMP_SIGNAL_9(24);
BusMuxIn-R1023 <= GDFX_TEMP_SIGNAL_9(23);
BusMuxIn-R1022 <= GDFX_TEMP_SIGNAL_9(22);
BusMuxIn-R1021 <= GDFX_TEMP_SIGNAL_9(21);
BusMuxIn-R1020 <= GDFX_TEMP_SIGNAL_9(20);
BusMuxIn-R1019 <= GDFX_TEMP_SIGNAL_9(19);
BusMuxIn-R1018 <= GDFX_TEMP_SIGNAL_9(18);
BusMuxIn-R1017 <= GDFX_TEMP_SIGNAL_9(17);
BusMuxIn-R1016 <= GDFX_TEMP_SIGNAL_9(16);
BusMuxIn-R1015 <= GDFX_TEMP_SIGNAL_9(15);
BusMuxIn-R1014 <= GDFX_TEMP_SIGNAL_9(14);
BusMuxIn-R1013 <= GDFX_TEMP_SIGNAL_9(13);
BusMuxIn-R1012 <= GDFX_TEMP_SIGNAL_9(12);
BusMuxIn-R1011 <= GDFX_TEMP_SIGNAL_9(11);
BusMuxIn-R1010 <= GDFX_TEMP_SIGNAL_9(10);
BusMuxIn-R109 <= GDFX_TEMP_SIGNAL_9(9);
BusMuxIn-R108 <= GDFX_TEMP_SIGNAL_9(8);
BusMuxIn-R107 <= GDFX_TEMP_SIGNAL_9(7);
BusMuxIn-R106 <= GDFX_TEMP_SIGNAL_9(6);
BusMuxIn-R105 <= GDFX_TEMP_SIGNAL_9(5);
BusMuxIn-R104 <= GDFX_TEMP_SIGNAL_9(4);
BusMuxIn-R103 <= GDFX_TEMP_SIGNAL_9(3);
BusMuxIn-R102 <= GDFX_TEMP_SIGNAL_9(2);
BusMuxIn-R101 <= GDFX_TEMP_SIGNAL_9(1);
BusMuxIn-R100 <= GDFX_TEMP_SIGNAL_9(0);

GDFX_TEMP_SIGNAL_6 <= (BusMuxIn-R131 & BusMuxIn-R130 & BusMuxIn-R129 & BusMuxIn-R128 & BusMuxIn-R127 & BusMuxIn-R126 & BusMuxIn-R125 & BusMuxIn-R124 & BusMuxIn-R123 & BusMuxIn-R122 & BusMuxIn-R121 & BusMuxIn-R120 & BusMuxIn-R119 & BusMuxIn-R118 & BusMuxIn-R117 & BusMuxIn-R116 & BusMuxIn-R115 & BusMuxIn-R114 & BusMuxIn-R113 & BusMuxIn-R112 & BusMuxIn-R111 & BusMuxIn-R110 & BusMuxIn-R19 & BusMuxIn-R18 & BusMuxIn-R17 & BusMuxIn-R16 & BusMuxIn-R15 & BusMuxIn-R14 & BusMuxIn-R13 & BusMuxIn-R12 & BusMuxIn-R11 & BusMuxIn-R10);
BusMuxIn-R131 <= GDFX_TEMP_SIGNAL_8(31);
BusMuxIn-R130 <= GDFX_TEMP_SIGNAL_8(30);
BusMuxIn-R129 <= GDFX_TEMP_SIGNAL_8(29);
BusMuxIn-R128 <= GDFX_TEMP_SIGNAL_8(28);
BusMuxIn-R127 <= GDFX_TEMP_SIGNAL_8(27);
BusMuxIn-R126 <= GDFX_TEMP_SIGNAL_8(26);
BusMuxIn-R125 <= GDFX_TEMP_SIGNAL_8(25);
BusMuxIn-R124 <= GDFX_TEMP_SIGNAL_8(24);
BusMuxIn-R123 <= GDFX_TEMP_SIGNAL_8(23);
BusMuxIn-R122 <= GDFX_TEMP_SIGNAL_8(22);
BusMuxIn-R121 <= GDFX_TEMP_SIGNAL_8(21);
BusMuxIn-R120 <= GDFX_TEMP_SIGNAL_8(20);
BusMuxIn-R119 <= GDFX_TEMP_SIGNAL_8(19);
BusMuxIn-R118 <= GDFX_TEMP_SIGNAL_8(18);
BusMuxIn-R117 <= GDFX_TEMP_SIGNAL_8(17);
BusMuxIn-R116 <= GDFX_TEMP_SIGNAL_8(16);
BusMuxIn-R115 <= GDFX_TEMP_SIGNAL_8(15);
BusMuxIn-R114 <= GDFX_TEMP_SIGNAL_8(14);
BusMuxIn-R113 <= GDFX_TEMP_SIGNAL_8(13);
BusMuxIn-R112 <= GDFX_TEMP_SIGNAL_8(12);
BusMuxIn-R111 <= GDFX_TEMP_SIGNAL_8(11);
BusMuxIn-R110 <= GDFX_TEMP_SIGNAL_8(10);
BusMuxIn-R19 <= GDFX_TEMP_SIGNAL_8(9);
BusMuxIn-R18 <= GDFX_TEMP_SIGNAL_8(8);
BusMuxIn-R17 <= GDFX_TEMP_SIGNAL_8(7);
BusMuxIn-R16 <= GDFX_TEMP_SIGNAL_8(6);
BusMuxIn-R15 <= GDFX_TEMP_SIGNAL_8(5);
BusMuxIn-R14 <= GDFX_TEMP_SIGNAL_8(4);
BusMuxIn-R13 <= GDFX_TEMP_SIGNAL_8(3);
BusMuxIn-R12 <= GDFX_TEMP_SIGNAL_8(2);
BusMuxIn-R11 <= GDFX_TEMP_SIGNAL_8(1);
BusMuxIn-R10 <= GDFX_TEMP_SIGNAL_8(0);

GDFX_TEMP_SIGNAL_7 <= (BusMuxIn-MDR31 & BusMuxIn-MDR30 & BusMuxIn-MDR29 & BusMuxIn-MDR28 & BusMuxIn-MDR27 & BusMuxIn-MDR26 & BusMuxIn-MDR25 & BusMuxIn-MDR24 & BusMuxIn-MDR23 & BusMuxIn-MDR22 & BusMuxIn-MDR21 & BusMuxIn-MDR20 & BusMuxIn-MDR19 & BusMuxIn-MDR18 & BusMuxIn-MDR17 & BusMuxIn-MDR16 & BusMuxIn-MDR15 & BusMuxIn-MDR14 & BusMuxIn-MDR13 & BusMuxIn-MDR12 & BusMuxIn-MDR11 & BusMuxIn-MDR10 & BusMuxIn-MDR9 & BusMuxIn-MDR8 & BusMuxIn-MDR7 & BusMuxIn-MDR6 & BusMuxIn-MDR5 & BusMuxIn-MDR4 & BusMuxIn-MDR3 & BusMuxIn-MDR2 & BusMuxIn-MDR1 & BusMuxIn-MDR0);


b2v_inst : lpm_encoder
PORT MAP(eq0 => R0out,
		 eq1 => R1out,
		 eq2 => R2out,
		 eq3 => R3out,
		 eq4 => R4out,
		 eq5 => R5out,
		 eq6 => R6out,
		 eq7 => R7out,
		 eq8 => R8out,
		 eq9 => R9out,
		 eq10 => R10out,
		 eq11 => R11out,
		 eq12 => R12out,
		 eq13 => R13out,
		 eq14 => R14out,
		 eq15 => R15out,
		 eq16 => HIout,
		 eq17 => LOout,
		 eq18 => Zhighout,
		 eq19 => Zlowout,
		 eq20 => PCout,
		 eq21 => MDRout,
		 eq22 => In_Portout,
		 eq23 => Cout,
		 data => muxSelect);


b2v_inst2 : lpm_mux0
PORT MAP(data0x => BusMuxIn-R0,
		 data10x => GDFX_TEMP_SIGNAL_0,
		 data11x => GDFX_TEMP_SIGNAL_1,
		 data12x => GDFX_TEMP_SIGNAL_2,
		 data13x => GDFX_TEMP_SIGNAL_3,
		 data14x => GDFX_TEMP_SIGNAL_4,
		 data15x => GDFX_TEMP_SIGNAL_5,
		 data16x => BusMuxIn-Hi,
		 data17x => BusMuxIn-Lo,
		 data18x => BusMuxIn-ZHi,
		 data19x => BusMuxIn-ZLo,
		 data1x => GDFX_TEMP_SIGNAL_6,
		 data20x => BusMuxIn-PC,
		 data21x => GDFX_TEMP_SIGNAL_7,
		 data22x => BusMuxIn-In_Port,
		 data23x => BusMuxIn-In_Port,
		 data2x => BusMuxIn-R2,
		 data3x => BusMuxIn-R3,
		 data4x => BusMuxIn-R4,
		 data5x => BusMuxIn-R5,
		 data6x => BusMuxIn-R6,
		 data7x => BusMuxIn-R7,
		 data8x => BusMuxIn-R8,
		 data9x => BusMuxIn-R9,
		 sel => muxSelect,
		 result => BusMuxOut);


b2v_MDR_Unit : mdr_unit
PORT MAP(MDR_IN_0 => BusMuxOut,
		 MDR_IN_1 => Mdatain);


b2v_REG0 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-R0);


b2v_REG1 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => GDFX_TEMP_SIGNAL_8);


b2v_REG10 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => GDFX_TEMP_SIGNAL_9);


b2v_REG11 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => GDFX_TEMP_SIGNAL_10);


b2v_REG12 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => GDFX_TEMP_SIGNAL_11);


b2v_REG13 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => GDFX_TEMP_SIGNAL_12);


b2v_REG14 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => GDFX_TEMP_SIGNAL_13);


b2v_REG15 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => GDFX_TEMP_SIGNAL_14);


b2v_REG2 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-R2);


b2v_REG3 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-R3);


b2v_REG4 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-R4);


b2v_REG5 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-R5);


b2v_REG6 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-R6);


b2v_REG7 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-R7);


b2v_REG8 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-R8);


b2v_REG9 : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-R9);


b2v_REGC : reg32
PORT MAP(D_IN => BusMuxOut);


b2v_REGHi : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-Hi);


b2v_REGIn_Port : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-In_Port);


b2v_REGLo : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-Lo);


b2v_REGPC : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-PC);


b2v_REGZHI : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-ZHi);


b2v_REGZLO : reg32
PORT MAP(D_IN => BusMuxOut,
		 D_OUT => BusMuxIn-ZLo);


BusMuxIn-R10 <= GDFX_TEMP_SIGNAL_8(0);
BusMuxIn-R100 <= GDFX_TEMP_SIGNAL_9(0);
BusMuxIn-R101 <= GDFX_TEMP_SIGNAL_9(1);
BusMuxIn-R1010 <= GDFX_TEMP_SIGNAL_9(10);
BusMuxIn-R1011 <= GDFX_TEMP_SIGNAL_9(11);
BusMuxIn-R1012 <= GDFX_TEMP_SIGNAL_9(12);
BusMuxIn-R1013 <= GDFX_TEMP_SIGNAL_9(13);
BusMuxIn-R1014 <= GDFX_TEMP_SIGNAL_9(14);
BusMuxIn-R1015 <= GDFX_TEMP_SIGNAL_9(15);
BusMuxIn-R1016 <= GDFX_TEMP_SIGNAL_9(16);
BusMuxIn-R1017 <= GDFX_TEMP_SIGNAL_9(17);
BusMuxIn-R1018 <= GDFX_TEMP_SIGNAL_9(18);
BusMuxIn-R1019 <= GDFX_TEMP_SIGNAL_9(19);
BusMuxIn-R102 <= GDFX_TEMP_SIGNAL_9(2);
BusMuxIn-R1020 <= GDFX_TEMP_SIGNAL_9(20);
BusMuxIn-R1021 <= GDFX_TEMP_SIGNAL_9(21);
BusMuxIn-R1022 <= GDFX_TEMP_SIGNAL_9(22);
BusMuxIn-R1023 <= GDFX_TEMP_SIGNAL_9(23);
BusMuxIn-R1024 <= GDFX_TEMP_SIGNAL_9(24);
BusMuxIn-R1025 <= GDFX_TEMP_SIGNAL_9(25);
BusMuxIn-R1026 <= GDFX_TEMP_SIGNAL_9(26);
BusMuxIn-R1027 <= GDFX_TEMP_SIGNAL_9(27);
BusMuxIn-R1028 <= GDFX_TEMP_SIGNAL_9(28);
BusMuxIn-R1029 <= GDFX_TEMP_SIGNAL_9(29);
BusMuxIn-R103 <= GDFX_TEMP_SIGNAL_9(3);
BusMuxIn-R1030 <= GDFX_TEMP_SIGNAL_9(30);
BusMuxIn-R1031 <= GDFX_TEMP_SIGNAL_9(31);
BusMuxIn-R104 <= GDFX_TEMP_SIGNAL_9(4);
BusMuxIn-R105 <= GDFX_TEMP_SIGNAL_9(5);
BusMuxIn-R106 <= GDFX_TEMP_SIGNAL_9(6);
BusMuxIn-R107 <= GDFX_TEMP_SIGNAL_9(7);
BusMuxIn-R108 <= GDFX_TEMP_SIGNAL_9(8);
BusMuxIn-R109 <= GDFX_TEMP_SIGNAL_9(9);
BusMuxIn-R11 <= GDFX_TEMP_SIGNAL_8(1);
BusMuxIn-R110 <= GDFX_TEMP_SIGNAL_10(0);
BusMuxIn-R110 <= GDFX_TEMP_SIGNAL_8(10);
BusMuxIn-R111 <= GDFX_TEMP_SIGNAL_10(1);
BusMuxIn-R111 <= GDFX_TEMP_SIGNAL_8(11);
BusMuxIn-R1110 <= GDFX_TEMP_SIGNAL_10(10);
BusMuxIn-R1111 <= GDFX_TEMP_SIGNAL_10(11);
BusMuxIn-R1112 <= GDFX_TEMP_SIGNAL_10(12);
BusMuxIn-R1113 <= GDFX_TEMP_SIGNAL_10(13);
BusMuxIn-R1114 <= GDFX_TEMP_SIGNAL_10(14);
BusMuxIn-R1115 <= GDFX_TEMP_SIGNAL_10(15);
BusMuxIn-R1116 <= GDFX_TEMP_SIGNAL_10(16);
BusMuxIn-R1117 <= GDFX_TEMP_SIGNAL_10(17);
BusMuxIn-R1118 <= GDFX_TEMP_SIGNAL_10(18);
BusMuxIn-R1119 <= GDFX_TEMP_SIGNAL_10(19);
BusMuxIn-R112 <= GDFX_TEMP_SIGNAL_10(2);
BusMuxIn-R112 <= GDFX_TEMP_SIGNAL_8(12);
BusMuxIn-R1120 <= GDFX_TEMP_SIGNAL_10(20);
BusMuxIn-R1121 <= GDFX_TEMP_SIGNAL_10(21);
BusMuxIn-R1122 <= GDFX_TEMP_SIGNAL_10(22);
BusMuxIn-R1123 <= GDFX_TEMP_SIGNAL_10(23);
BusMuxIn-R1124 <= GDFX_TEMP_SIGNAL_10(24);
BusMuxIn-R1125 <= GDFX_TEMP_SIGNAL_10(25);
BusMuxIn-R1126 <= GDFX_TEMP_SIGNAL_10(26);
BusMuxIn-R1127 <= GDFX_TEMP_SIGNAL_10(27);
BusMuxIn-R1128 <= GDFX_TEMP_SIGNAL_10(28);
BusMuxIn-R1129 <= GDFX_TEMP_SIGNAL_10(29);
BusMuxIn-R113 <= GDFX_TEMP_SIGNAL_10(3);
BusMuxIn-R113 <= GDFX_TEMP_SIGNAL_8(13);
BusMuxIn-R1130 <= GDFX_TEMP_SIGNAL_10(30);
BusMuxIn-R1131 <= GDFX_TEMP_SIGNAL_10(31);
BusMuxIn-R114 <= GDFX_TEMP_SIGNAL_10(4);
BusMuxIn-R114 <= GDFX_TEMP_SIGNAL_8(14);
BusMuxIn-R115 <= GDFX_TEMP_SIGNAL_10(5);
BusMuxIn-R115 <= GDFX_TEMP_SIGNAL_8(15);
BusMuxIn-R116 <= GDFX_TEMP_SIGNAL_10(6);
BusMuxIn-R116 <= GDFX_TEMP_SIGNAL_8(16);
BusMuxIn-R117 <= GDFX_TEMP_SIGNAL_10(7);
BusMuxIn-R117 <= GDFX_TEMP_SIGNAL_8(17);
BusMuxIn-R118 <= GDFX_TEMP_SIGNAL_10(8);
BusMuxIn-R118 <= GDFX_TEMP_SIGNAL_8(18);
BusMuxIn-R119 <= GDFX_TEMP_SIGNAL_10(9);
BusMuxIn-R119 <= GDFX_TEMP_SIGNAL_8(19);
BusMuxIn-R12 <= GDFX_TEMP_SIGNAL_8(2);
BusMuxIn-R120 <= GDFX_TEMP_SIGNAL_8(20);
BusMuxIn-R120 <= GDFX_TEMP_SIGNAL_11(0);
BusMuxIn-R121 <= GDFX_TEMP_SIGNAL_8(21);
BusMuxIn-R121 <= GDFX_TEMP_SIGNAL_11(1);
BusMuxIn-R1210 <= GDFX_TEMP_SIGNAL_11(10);
BusMuxIn-R1211 <= GDFX_TEMP_SIGNAL_11(11);
BusMuxIn-R1212 <= GDFX_TEMP_SIGNAL_11(12);
BusMuxIn-R1213 <= GDFX_TEMP_SIGNAL_11(13);
BusMuxIn-R1214 <= GDFX_TEMP_SIGNAL_11(14);
BusMuxIn-R1215 <= GDFX_TEMP_SIGNAL_11(15);
BusMuxIn-R1216 <= GDFX_TEMP_SIGNAL_11(16);
BusMuxIn-R1217 <= GDFX_TEMP_SIGNAL_11(17);
BusMuxIn-R1218 <= GDFX_TEMP_SIGNAL_11(18);
BusMuxIn-R1219 <= GDFX_TEMP_SIGNAL_11(19);
BusMuxIn-R122 <= GDFX_TEMP_SIGNAL_8(22);
BusMuxIn-R122 <= GDFX_TEMP_SIGNAL_11(2);
BusMuxIn-R1220 <= GDFX_TEMP_SIGNAL_11(20);
BusMuxIn-R1221 <= GDFX_TEMP_SIGNAL_11(21);
BusMuxIn-R1222 <= GDFX_TEMP_SIGNAL_11(22);
BusMuxIn-R1223 <= GDFX_TEMP_SIGNAL_11(23);
BusMuxIn-R1224 <= GDFX_TEMP_SIGNAL_11(24);
BusMuxIn-R1225 <= GDFX_TEMP_SIGNAL_11(25);
BusMuxIn-R1226 <= GDFX_TEMP_SIGNAL_11(26);
BusMuxIn-R1227 <= GDFX_TEMP_SIGNAL_11(27);
BusMuxIn-R1228 <= GDFX_TEMP_SIGNAL_11(28);
BusMuxIn-R1229 <= GDFX_TEMP_SIGNAL_11(29);
BusMuxIn-R123 <= GDFX_TEMP_SIGNAL_8(23);
BusMuxIn-R123 <= GDFX_TEMP_SIGNAL_11(3);
BusMuxIn-R1230 <= GDFX_TEMP_SIGNAL_11(30);
BusMuxIn-R1231 <= GDFX_TEMP_SIGNAL_11(31);
BusMuxIn-R124 <= GDFX_TEMP_SIGNAL_8(24);
BusMuxIn-R124 <= GDFX_TEMP_SIGNAL_11(4);
BusMuxIn-R125 <= GDFX_TEMP_SIGNAL_8(25);
BusMuxIn-R125 <= GDFX_TEMP_SIGNAL_11(5);
BusMuxIn-R126 <= GDFX_TEMP_SIGNAL_8(26);
BusMuxIn-R126 <= GDFX_TEMP_SIGNAL_11(6);
BusMuxIn-R127 <= GDFX_TEMP_SIGNAL_8(27);
BusMuxIn-R127 <= GDFX_TEMP_SIGNAL_11(7);
BusMuxIn-R128 <= GDFX_TEMP_SIGNAL_8(28);
BusMuxIn-R128 <= GDFX_TEMP_SIGNAL_11(8);
BusMuxIn-R129 <= GDFX_TEMP_SIGNAL_8(29);
BusMuxIn-R129 <= GDFX_TEMP_SIGNAL_11(9);
BusMuxIn-R13 <= GDFX_TEMP_SIGNAL_8(3);
BusMuxIn-R130 <= GDFX_TEMP_SIGNAL_8(30);
BusMuxIn-R130 <= GDFX_TEMP_SIGNAL_12(0);
BusMuxIn-R131 <= GDFX_TEMP_SIGNAL_8(31);
BusMuxIn-R131 <= GDFX_TEMP_SIGNAL_12(1);
BusMuxIn-R1310 <= GDFX_TEMP_SIGNAL_12(10);
BusMuxIn-R1311 <= GDFX_TEMP_SIGNAL_12(11);
BusMuxIn-R1312 <= GDFX_TEMP_SIGNAL_12(12);
BusMuxIn-R1313 <= GDFX_TEMP_SIGNAL_12(13);
BusMuxIn-R1314 <= GDFX_TEMP_SIGNAL_12(14);
BusMuxIn-R1315 <= GDFX_TEMP_SIGNAL_12(15);
BusMuxIn-R1316 <= GDFX_TEMP_SIGNAL_12(16);
BusMuxIn-R1317 <= GDFX_TEMP_SIGNAL_12(17);
BusMuxIn-R1318 <= GDFX_TEMP_SIGNAL_12(18);
BusMuxIn-R1319 <= GDFX_TEMP_SIGNAL_12(19);
BusMuxIn-R132 <= GDFX_TEMP_SIGNAL_12(2);
BusMuxIn-R1320 <= GDFX_TEMP_SIGNAL_12(20);
BusMuxIn-R1321 <= GDFX_TEMP_SIGNAL_12(21);
BusMuxIn-R1322 <= GDFX_TEMP_SIGNAL_12(22);
BusMuxIn-R1323 <= GDFX_TEMP_SIGNAL_12(23);
BusMuxIn-R1324 <= GDFX_TEMP_SIGNAL_12(24);
BusMuxIn-R1325 <= GDFX_TEMP_SIGNAL_12(25);
BusMuxIn-R1326 <= GDFX_TEMP_SIGNAL_12(26);
BusMuxIn-R1327 <= GDFX_TEMP_SIGNAL_12(27);
BusMuxIn-R1328 <= GDFX_TEMP_SIGNAL_12(28);
BusMuxIn-R1329 <= GDFX_TEMP_SIGNAL_12(29);
BusMuxIn-R133 <= GDFX_TEMP_SIGNAL_12(3);
BusMuxIn-R1330 <= GDFX_TEMP_SIGNAL_12(30);
BusMuxIn-R1331 <= GDFX_TEMP_SIGNAL_12(31);
BusMuxIn-R134 <= GDFX_TEMP_SIGNAL_12(4);
BusMuxIn-R135 <= GDFX_TEMP_SIGNAL_12(5);
BusMuxIn-R136 <= GDFX_TEMP_SIGNAL_12(6);
BusMuxIn-R137 <= GDFX_TEMP_SIGNAL_12(7);
BusMuxIn-R138 <= GDFX_TEMP_SIGNAL_12(8);
BusMuxIn-R139 <= GDFX_TEMP_SIGNAL_12(9);
BusMuxIn-R14 <= GDFX_TEMP_SIGNAL_8(4);
BusMuxIn-R140 <= GDFX_TEMP_SIGNAL_13(0);
BusMuxIn-R141 <= GDFX_TEMP_SIGNAL_13(1);
BusMuxIn-R1410 <= GDFX_TEMP_SIGNAL_13(10);
BusMuxIn-R1411 <= GDFX_TEMP_SIGNAL_13(11);
BusMuxIn-R1412 <= GDFX_TEMP_SIGNAL_13(12);
BusMuxIn-R1413 <= GDFX_TEMP_SIGNAL_13(13);
BusMuxIn-R1414 <= GDFX_TEMP_SIGNAL_13(14);
BusMuxIn-R1415 <= GDFX_TEMP_SIGNAL_13(15);
BusMuxIn-R1416 <= GDFX_TEMP_SIGNAL_13(16);
BusMuxIn-R1417 <= GDFX_TEMP_SIGNAL_13(17);
BusMuxIn-R1418 <= GDFX_TEMP_SIGNAL_13(18);
BusMuxIn-R1419 <= GDFX_TEMP_SIGNAL_13(19);
BusMuxIn-R142 <= GDFX_TEMP_SIGNAL_13(2);
BusMuxIn-R1420 <= GDFX_TEMP_SIGNAL_13(20);
BusMuxIn-R1421 <= GDFX_TEMP_SIGNAL_13(21);
BusMuxIn-R1422 <= GDFX_TEMP_SIGNAL_13(22);
BusMuxIn-R1423 <= GDFX_TEMP_SIGNAL_13(23);
BusMuxIn-R1424 <= GDFX_TEMP_SIGNAL_13(24);
BusMuxIn-R1425 <= GDFX_TEMP_SIGNAL_13(25);
BusMuxIn-R1426 <= GDFX_TEMP_SIGNAL_13(26);
BusMuxIn-R1427 <= GDFX_TEMP_SIGNAL_13(27);
BusMuxIn-R1428 <= GDFX_TEMP_SIGNAL_13(28);
BusMuxIn-R1429 <= GDFX_TEMP_SIGNAL_13(29);
BusMuxIn-R143 <= GDFX_TEMP_SIGNAL_13(3);
BusMuxIn-R1430 <= GDFX_TEMP_SIGNAL_13(30);
BusMuxIn-R1431 <= GDFX_TEMP_SIGNAL_13(31);
BusMuxIn-R144 <= GDFX_TEMP_SIGNAL_13(4);
BusMuxIn-R145 <= GDFX_TEMP_SIGNAL_13(5);
BusMuxIn-R146 <= GDFX_TEMP_SIGNAL_13(6);
BusMuxIn-R147 <= GDFX_TEMP_SIGNAL_13(7);
BusMuxIn-R148 <= GDFX_TEMP_SIGNAL_13(8);
BusMuxIn-R149 <= GDFX_TEMP_SIGNAL_13(9);
BusMuxIn-R15 <= GDFX_TEMP_SIGNAL_8(5);
BusMuxIn-R150 <= GDFX_TEMP_SIGNAL_14(0);
BusMuxIn-R151 <= GDFX_TEMP_SIGNAL_14(1);
BusMuxIn-R1510 <= GDFX_TEMP_SIGNAL_14(10);
BusMuxIn-R1511 <= GDFX_TEMP_SIGNAL_14(11);
BusMuxIn-R1512 <= GDFX_TEMP_SIGNAL_14(12);
BusMuxIn-R1513 <= GDFX_TEMP_SIGNAL_14(13);
BusMuxIn-R1514 <= GDFX_TEMP_SIGNAL_14(14);
BusMuxIn-R1515 <= GDFX_TEMP_SIGNAL_14(15);
BusMuxIn-R1516 <= GDFX_TEMP_SIGNAL_14(16);
BusMuxIn-R1517 <= GDFX_TEMP_SIGNAL_14(17);
BusMuxIn-R1518 <= GDFX_TEMP_SIGNAL_14(18);
BusMuxIn-R1519 <= GDFX_TEMP_SIGNAL_14(19);
BusMuxIn-R152 <= GDFX_TEMP_SIGNAL_14(2);
BusMuxIn-R1520 <= GDFX_TEMP_SIGNAL_14(20);
BusMuxIn-R1521 <= GDFX_TEMP_SIGNAL_14(21);
BusMuxIn-R1522 <= GDFX_TEMP_SIGNAL_14(22);
BusMuxIn-R1523 <= GDFX_TEMP_SIGNAL_14(23);
BusMuxIn-R1524 <= GDFX_TEMP_SIGNAL_14(24);
BusMuxIn-R1525 <= GDFX_TEMP_SIGNAL_14(25);
BusMuxIn-R1526 <= GDFX_TEMP_SIGNAL_14(26);
BusMuxIn-R1527 <= GDFX_TEMP_SIGNAL_14(27);
BusMuxIn-R1528 <= GDFX_TEMP_SIGNAL_14(28);
BusMuxIn-R1529 <= GDFX_TEMP_SIGNAL_14(29);
BusMuxIn-R153 <= GDFX_TEMP_SIGNAL_14(3);
BusMuxIn-R1530 <= GDFX_TEMP_SIGNAL_14(30);
BusMuxIn-R1531 <= GDFX_TEMP_SIGNAL_14(31);
BusMuxIn-R154 <= GDFX_TEMP_SIGNAL_14(4);
BusMuxIn-R155 <= GDFX_TEMP_SIGNAL_14(5);
BusMuxIn-R156 <= GDFX_TEMP_SIGNAL_14(6);
BusMuxIn-R157 <= GDFX_TEMP_SIGNAL_14(7);
BusMuxIn-R158 <= GDFX_TEMP_SIGNAL_14(8);
BusMuxIn-R159 <= GDFX_TEMP_SIGNAL_14(9);
BusMuxIn-R16 <= GDFX_TEMP_SIGNAL_8(6);
BusMuxIn-R17 <= GDFX_TEMP_SIGNAL_8(7);
BusMuxIn-R18 <= GDFX_TEMP_SIGNAL_8(8);
BusMuxIn-R19 <= GDFX_TEMP_SIGNAL_8(9);
END bdf_type;