package Common is

type State IS (Reset_state, 
							fetch0, 
							fetch1, 
							fetch2,
							addImmediate3,
							addImmediate4,
							addImmediate5,
							addImmediate6,
							zero,
							add3, 
							add4, 
							add5, 
							add6, 
							load3, 
							load4, 
							load5, 
							load6, 
							load7, 
							loadImmediate3, 
							loadImmediate4, 
							loadImmediate5,
							loadRelative3,
							loadRelative4,
							loadRelative5,
							loadRelative6,
							andImmediate3,
							andImmediate4,
							andImmediate5,
							sub3,
							sub4,
							sub5,
							negate3,
							negate4,
							negate5,
							not3,
							not4,
							not5,
							shr3,
							shr4,
							shr5,
							shl3,
							shl4,
							shl5,
							ror3,
							ror4,
							ror5,
							rol3,
							rol4,
							rol5,
							or3,
							or4,
							or5,
							and3,
							and4,
							and5,
							multiply3,
							multiply4,
							multiply5,
							multiply6,
							divide3,
							divide4,
							divide5,
							divide6,
							mfhi3,
							mflo3,
							jal3,
							jal4,
							jal5,
							jr3,
							orImmediate3,
							orImmediate4,
							orImmediate5,
							storeRelative3,
							storeRelative4,
							storeRelative5,
							storeRelative6,
							storeRelative7,
							store3,
							store4,
							store5,
							store6,
							store7,
							out3,
							in3,
							in4,
							brzr3,
							brzr4,
							brnz3,
							brnz4,
							halt,
							nop
							);

end Common;
